* AC Analysis Script
* Load the SPICE file
source basic_circuit.spice
* Run AC analysis
ac
* Print AC results
print all
* End of script
.end

