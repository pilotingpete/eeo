* DC Analysis Script
* Load the SPICE file
source basic_circuit.spice
* Run DC analysis
op
* Print DC operating point
print all
* End of script
.end
