** Profile: "SCHEMATIC1-PMsweep"  [ c:\cds_spb_home\cdssetup\projects\pm-sim1\pm-sim1-PSpiceFiles\SCHEMATIC1\PMsweep.sim ] 

** Creating circuit file "PMsweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/eeo/eeo-311/simulation/s-1/ese311models.lib" 
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 1 .01 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
