* First-Order Low-Pass Filter

* Input voltage source
Vin N1 0 AC 1V SIN(0 1V 10kHz)  ; 1V amplitude AC voltage source at node 1 (input)

* Define the components
R1 N1 N2 1k  ; 1.0k ohm resistor
C1 N2 0 4.7n ; 4.7 nF capacitor

* AC analysis
.ac dec 10 1 100k  ; AC sweep 

* Node N2: Output Node

* Analysis
.control
  run
  plot mag(N2)  ; Bode plot of the magnitude of Vout
  plot phase(N2)  ; Bode plot of the phase of Vout
.endc

.end
